library verilog;
use verilog.vl_types.all;
entity projetoProcessador is
    generic(
        T0              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        T1              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        T2              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        T3              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        T4              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        T5              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        mv              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        mvt             : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        add             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        sub             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        load            : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        store           : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        \_and\          : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        b_cond          : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        shift           : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        \_R0\           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        \_R1\           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        \_R2\           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        \_R3\           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        \_R4\           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        \_R5\           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        \_R6\           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        \_PC\           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        \_G\            : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        \_IR8_IR8_0\    : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        \_IR7_0_0\      : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        \_DIN\          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1)
    );
    port(
        Resetn          : in     vl_logic;
        Clock           : in     vl_logic;
        Run             : in     vl_logic;
        Done            : out    vl_logic;
        reg0            : out    vl_logic_vector(15 downto 0);
        reg1            : out    vl_logic_vector(15 downto 0);
        reg2            : out    vl_logic_vector(15 downto 0);
        reg3            : out    vl_logic_vector(15 downto 0);
        reg4            : out    vl_logic_vector(15 downto 0);
        reg5            : out    vl_logic_vector(15 downto 0);
        reg6            : out    vl_logic_vector(15 downto 0);
        regPC           : out    vl_logic_vector(15 downto 0);
        Instr           : out    vl_logic_vector(15 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of T0 : constant is 1;
    attribute mti_svvh_generic_type of T1 : constant is 1;
    attribute mti_svvh_generic_type of T2 : constant is 1;
    attribute mti_svvh_generic_type of T3 : constant is 1;
    attribute mti_svvh_generic_type of T4 : constant is 1;
    attribute mti_svvh_generic_type of T5 : constant is 1;
    attribute mti_svvh_generic_type of mv : constant is 1;
    attribute mti_svvh_generic_type of mvt : constant is 1;
    attribute mti_svvh_generic_type of add : constant is 1;
    attribute mti_svvh_generic_type of sub : constant is 1;
    attribute mti_svvh_generic_type of load : constant is 1;
    attribute mti_svvh_generic_type of store : constant is 1;
    attribute mti_svvh_generic_type of \_and\ : constant is 1;
    attribute mti_svvh_generic_type of b_cond : constant is 1;
    attribute mti_svvh_generic_type of shift : constant is 1;
    attribute mti_svvh_generic_type of \_R0\ : constant is 1;
    attribute mti_svvh_generic_type of \_R1\ : constant is 1;
    attribute mti_svvh_generic_type of \_R2\ : constant is 1;
    attribute mti_svvh_generic_type of \_R3\ : constant is 1;
    attribute mti_svvh_generic_type of \_R4\ : constant is 1;
    attribute mti_svvh_generic_type of \_R5\ : constant is 1;
    attribute mti_svvh_generic_type of \_R6\ : constant is 1;
    attribute mti_svvh_generic_type of \_PC\ : constant is 1;
    attribute mti_svvh_generic_type of \_G\ : constant is 1;
    attribute mti_svvh_generic_type of \_IR8_IR8_0\ : constant is 1;
    attribute mti_svvh_generic_type of \_IR7_0_0\ : constant is 1;
    attribute mti_svvh_generic_type of \_DIN\ : constant is 1;
end projetoProcessador;
