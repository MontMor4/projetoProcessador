library verilog;
use verilog.vl_types.all;
entity projetoProcessador_tb is
end projetoProcessador_tb;
